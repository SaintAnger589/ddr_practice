module command_top (

);


//signal interface

//arbiter

//multiplexer

//shift registers



endmodule